** Profile: "SCHEMATIC1-test"  [ H:\Uni Stuff\Year 3\Project\Pspice\test AD549\test AD549-PSpiceFiles\SCHEMATIC1\test.sim ] 

** Creating circuit file "test.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "H:/Uni Stuff/Year 3/Project/Pspice/models/opa124_pspice_aio/opa124.lib" 
.LIB "H:/Uni Stuff/Year 3/Project/Pspice/models/ad549/ad549.lib" 
* From [PSPICE NETLIST] section of H:\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN I_I1 0 100p 0.001p 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
